module TRANS(
    getinst_inst_i,
    trans_instruct_o,
    dmem_rs1_o,
    dmem_rs2_o,
    clk_i,
    rst_n_i
)

wire clk_i;
wire rst_n_i;